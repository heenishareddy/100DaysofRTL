`timescale 1ns / 1ps

module fulladdertb;
  reg a, b, cin;
  wire sout, cout;

  fulladder dut(a, b, cin, sout, cout);

  initial begin
    clk = 0;
    a = 0; b = 0; cin = 0;
    #10;
    a = 0; b = 0; cin = 1;
    #10;
    a = 0; b = 1; cin = 0;
    #10;
    a = 0; b = 1; cin = 1;
    #10;
    a = 1; b = 0; cin = 0;
    #10;
    a = 1; b = 0; cin = 1;
    #10;
    a = 1; b = 1; cin = 0;
    #10;
    a = 1; b = 1; cin = 1;
    #10;
    
  end